//=============================================================
// SHA-256 Initial Hash Values (FIPS 180-4, Section 5.3.3)
//=============================================================

`define H1_INIT 32'h6a09e667
`define H2_INIT 32'hbb67ae85
`define H3_INIT 32'h3c6ef372
`define H4_INIT 32'ha54ff53a
`define H5_INIT 32'h510e527f
`define H6_INIT 32'h9b05688c
`define H7_INIT 32'h1f83d9ab
`define H8_INIT 32'h5be0cd19

